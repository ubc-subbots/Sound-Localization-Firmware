//=================================
// Toggle on and off the desired properties for self checking

// `define NO_TIMING