//=================================
// Toggle on and off the desired properties for self checking

// ADC property checks
`define VALID_CHANNEL // check that ADC channel never goes above 5