// Analog waveform signal generation

