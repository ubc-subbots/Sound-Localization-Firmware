// Write Access Timing
`define tCSWR
`define tWRL
`define tWRH
`define tWRCS
`define tSUDI
`define tHDI


// Read Access Timing
`define tCONV 1330
`define tDCVB 25
`define tCVL  20
`define tRDL  20
`define tPDDO 15